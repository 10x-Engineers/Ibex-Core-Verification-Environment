// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

package mem_model_pkg;

  import uvm_pkg::*;

  `include "uvm_macros.svh"
  `include "verif/mem_model.sv"

endpackage
